//------------------
//  hogehoge
//------------------
module hogehoge(
);
endmodule


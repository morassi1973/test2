module newfile(
);
endmodule

